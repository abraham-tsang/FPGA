library ieee;
use ieee.std_logic_1164.all;

entity Subtractor is
    port (a, b : in std_logic_vector(3 downto 0); s : out std_logic_vector(3 downto 0));
end Subtractor;

architecture basic of Subtractor is
begin
    
end architecture basic;
